`timescale 1ns / 1ps

module ROM (
    input  logic [31:0] addr,
    output logic [31:0] data
);
    logic [31:0] rom[0:2**8-1];

    // 0   1    2   3   4   5    6    7     8   9
    // 10, 11, 12, 13, 14, -10, -11, -12, -13, -14

    initial begin
        // $readmemh("code.mem", rom);

        //rom[x]=32'b fucn7 _ rs2 _ rs1 _f3 _ rd  _ op // R-Type
        rom[0] = 32'b0000000_00001_00010_000_01010_0110011;  // add x10, x2, x1
        rom[1] = 32'b0100000_00001_00100_000_01011_0110011;  // sub x11, x4, x1
        rom[2] = 32'b0000000_00000_00011_111_01100_0110011;  // and x12, x3, x0
        rom[3] = 32'b0000000_00000_00011_110_01101_0110011;  // or  x13, x3, x0
        rom[4] = 32'b0100000_01011_00110_101_01110_0110011;  // sra x14, x6, x11
        rom[5] = 32'b0100000_01011_00111_101_01111_0110011;  // sra x15, x7, x11
        // rom[6] = 32'b0100000_01111_10000_101_10000_0110011;  // sra x16, x16, x15
        rom[6] = 32'b0000000_01011_01000_001_10000_0110011;  // sll x16, x8, x11
        rom[7] = 32'b0000000_01011_01000_101_10001_0110011;  // srl x17, x8, x11
        rom[8] = 32'b0000000_00000_00011_100_10010_0110011;  // bitxor x18, x3, x0
        rom[9] = 32'b0000000_00001_01001_010_10011_0110011;  // slt x19, x9, x1 (-14 < 14) 1
        // rom[10] = 32'b0000000_00000_01010_010_10101_0110011; // slt x21, x10, x0 (10 < 0) 0
        rom[10] = 32'b0000000_00001_01001_011_10100_0110011; // sltu x20, x9, x1 (-14 < 14) 0
        rom[12] = 32'b0000000_00000_10000_011_10101_0110011; // sltu x21, x16, x0 (unsigned(-10) < 0) 0
        rom[13] = 32'b0100000_00011_00001_000_01011_0110011;  // sub x11, x1, x3
        //rom[x]=32'b imm12      _ rs1 _f3 _ rd  _ op // I-Type  rd, rs1, imm
        rom[11] = 32'b0000000_00001_00001_000_10101_0010011;  // addi x21, x1, 1 
        rom[12] = 32'b0000000_00100_00011_111_10110_0010011;  // andi x22, x3, 4 
        rom[13] = 32'b0000000_00001_00011_110_10111_0010011;  // ori x23, x3, 1
        rom[14] = 32'b0000000_00011_01000_001_11000_0010011; // slli x24, x8, 3 // 2b00001011 << 3      1011000
        rom[15] = 32'b0000000_00100_01000_101_11001_0010011; // srli, x25, x8, 4 => regfile[13] = regfile[2] >> 4
        rom[16] = 32'b0100000_00011_00110_101_11010_0010011; // srai, x26, x6, 4 => regfile[20] = regfile[16] >>> 4
        rom[17] = 32'b0000000_00100_01001_010_11011_0010011; // slti, x27, x9, 4 => regfile[14] = regfile[3] < 4    1
        rom[18] = 32'b0000000_00100_01001_011_11100_0010011; // sltiu, x28, x9, 4 => regfile[15] = regfile[3] < 4  0
        rom[19] = 32'b0000000_00001_00011_100_11101_0010011; // xori, x29, x3, 1 => regfile[31] = regfile[3] ^ (11100000)
        // LU - Type                                               rd, imm
        rom[20] = 32'b00000000000000000001_11110_0110111;  // lui x30, 1 <<12
        // AU - Type                                                 rd, imm
        rom[21] = 32'b00000000000000000001_11111_0010111;  // auipc x31, 1   regfile[0] = pc+(1<<12) 'O'
        //rom[x]=32'b imm7  _ rs2 _ rs1 _f3 _ imm5_ op // S-Type    rs2, imm(rs1)
        rom[22] = 32'b0000000_00110_00000_010_01000_0100011;  // sw x6, 8(x0)
        rom[23] = 32'b0000000_00101_00100_110_01100_1100011;  // BLTU x4, x5 , 12
        rom[26] = 32'b0000000_00110_00000_000_00000_0100011; // sb x6, 0(x0) = rs1 + imm  ram[(0 + 0)>>2] = regfile[16]
        rom[27] = 32'b0000000_00100_00101_111_01100_1100011;  // BGEU x5, x4, 12
        rom[30] = 32'b0000000_00110_00000_001_00100_0100011; // sh x6, 4(x0) = rs1 + imm  ram[(0 + 4)>>2] = regfile[17]
        // // //rom[x]=32'b imm12      _ rs1 _f3 _ rd  _ op // L-Type  rd, imm(rs1)
        rom[31] = 32'b0000000_01000_00000_010_01010_0000011;// lw x10, 8(x0)    regfile[10] = ram[(0+8)/4]
        rom[32] = 32'b0000000_00010_00010_000_01100_1100011;  // beq x2, x2, 12
        rom[35] = 32'b0000000_00000_00000_000_01011_0000011; // lb, x11, 0(x0) => regfile[11] = ram[(0 + 0)>>2]
        rom[36] = 32'b0000000_00101_00110_001_01100_1100011;  // BNE  x5, x6, 12
        rom[39] = 32'b0000000_00100_00000_001_01101_0000011; // lh, x13, 4(x0) => regfile[13] = ram[(0 + 4)>>2]
        rom[40] = 32'b0000000_00100_00011_100_01100_1100011;  // BLT  x3, x4, 12
        rom[43] = 32'b0000000_00000_00000_100_01100_0000011; // lbu, x12, 0(x0) => regfile[12] = ram[(0 + 0)>>2]
        rom[44] = 32'b0000000_01001_01000_101_01100_1100011;  // BGE  x8, x9, 12
        rom[47] = 32'b0000000_00100_00000_101_01110_0000011; // lhu, x14, 4(x0) => regfile[14] = ram[(0 + 4)>>2]
        rom[48] = 32'b0000000_00110_00000_000_00001_0100011; // sb x6, 1(x0) = rs1 + imm  ram[(0 + 1)>>2] = regfile[16]
        rom[49] = 32'b0000000_00110_00000_000_00010_0100011; // sb x6, 2(x0) = rs1 + imm  ram[(0 + 2)>>2] = regfile[16]
        rom[50] = 32'b0000000_00110_00000_000_00011_0100011; // sb x6, 3(x0) = rs1 + imm  ram[(0 + 3)>>2] = regfile[16]
        // rom[51] = 32'b0000000_00110_00000_001_00101_0100011; // sh x6, 5(x0) = rs1 + imm  ram[(0 + 0)>>2] = regfile[16] -> 의도적 불량 명령어
        rom[51] = 32'b0000000_00110_00000_001_00110_0100011; // sh x6, 6(x0) = rs1 + imm  ram[(0 + 6)>>2] = regfile[16]
        rom[52] = 32'b0000000_00100_00000_001_01101_0000011; // lh, x13, 4(x0) => regfile[13] = ram[(0 + 4)>>2]
        rom[53] = 32'b0000000_00000_00000_100_01100_0000011; // lbu, x12, 0(x0) => regfile[12] = ram[(0 + 0)>>2]
        rom[54] = 32'b0000000_00110_00000_001_01101_0100011; // sh x6, 13(x0) = rs1 + imm  ram[(0 + 13)>>2] = regfile[6]
        rom[55] = 32'b0000000_00110_00000_001_01111_0100011; // sh x6, 15(x0) = rs1 + imm  ram[(0 + 15)>>2] = regfile[6]  // 저장 안함
        rom[56] = 32'b0000000_00101_00000_000_01111_0000011; // lb, x15, 5(x0) => regfile[11] = ram[(0 + 5)>>2]
        rom[57] = 32'b0000000_00110_00000_000_10000_0000011; // lb, x16, 6(x0) => regfile[11] = ram[(0 + 6)>>2]
        rom[58] = 32'b0000000_00111_00000_000_10001_0000011; // lb, x17, 7(x0) => regfile[11] = ram[(0 + 7)>>2]
        rom[59] = 32'b0000000_00101_00000_100_10010_0000011; // lbu, x18, 5(x0) => regfile[12] = ram[(0 + 5)>>2]
        rom[60] = 32'b0000000_00110_00000_100_10011_0000011; // lbu, x19, 6(x0) => regfile[12] = ram[(0 + 6)>>2]
        rom[61] = 32'b0000000_00111_00000_100_10100_0000011; // lbu, x20, 7(x0) => regfile[12] = ram[(0 + 7)>>2]
        rom[62] = 32'b0000000_01001_00000_001_10101_0000011; // lh, x21, 9(x0) => regfile[13] = ram[(0 + 9)>>2]
        rom[63] = 32'b0000000_01010_00000_001_10110_0000011; // lh, x22, 10(x0) => regfile[13] = ram[(0 + 10)>>2]
        rom[64] = 32'b0000000_01011_00000_001_10111_0000011; // lh, x23, 11(x0) => regfile[13] = ram[(0 + 11)>>2] // 안 가져옴
        rom[65] = 32'b0000000_01001_00000_101_11000_0000011; // lhu, x24, 9(x0) => regfile[13] = ram[(0 + 9)>>2]
        rom[66] = 32'b0000000_01010_00000_101_11001_0000011; // lhu, x25, 10(x0) => regfile[13] = ram[(0 + 10)>>2]
        rom[67] = 32'b0000000_01011_00000_101_11010_0000011; // lhu, x26, 11(x0) => regfile[13] = ram[(0 + 11)>>2] // 안 가져옴

        // rom[0] = 32'b0_0000000100_0_00000000_00001_1101111; // J
        // rom[2] = 32'b000000001000_00001_000_00010_1100111; // JA

        // rom[0] = 32'b0000000_00010_00010_000_01100_1100011;  // beq x2, x2, 12
        // rom[3] = 32'b0000000_00101_00110_001_01100_1100011;  // BNE  x5, x6, 12
        // rom[6] = 32'b0000000_00100_00011_100_01100_1100011;  // BLT  x3, x4, 12
        // rom[9] = 32'b0000000_01001_01000_101_01100_1100011;  // BGE  x8, x9, 12
        // rom[12] = 32'b0000000_00101_00100_110_01100_1100011;  // BLTU x4, x5 , 12
        // rom[15] = 32'b0000000_00100_00101_111_01100_1100011;  // BGEU x5, x4, 12
        // rom[6] = 
        // rom[7] =  // lhu, x14, 4(x0) => regfile[14] = ram[(0 + 4)>>2]
        // rom[8] = 32'b0000000_00001_00011_100_11101_0010011;
        // rom[9] = 
        // rom[10]= 
    end

    assign data = rom[addr[31:2]];
endmodule
