`timescale 1ns / 1ps

module CPU_RV32I (
    input  logic        clk,
    input  logic        reset,
    input  logic [31:0] instrCode,
    output logic [31:0] instrMemAddr,
    output logic        busWe,
    output logic [31:0] busAddr,
    output logic [31:0] busWData,
    input  logic [31:0] busRData,
    output logic [ 3:0] wstrb,
    output logic        st_misaligned
);
    logic       regFileWe;
    logic [3:0] aluControl;
    logic       aluSrcMuxSel;
    logic [2:0] RFWDSrcMuxSel;
    logic [2:0] LoadSizeMuxSel;
    logic [1:0] StoreSizeMuxSel;
    logic       branch;
    logic       jal;
    logic       jalr;
    logic       PCEn;


    ControlUnit U_ControlUnit (.*);
    DataPath U_DataPath (.*);
endmodule
